module phy
( 
 input ref_clk,
 input [1:0] tx_data,
 input tx_en,
 output [1:0] rx_data,
 output crs_dv,
 output rx_err
);
endmodule
